../../src/util/edge_detector.sv