../../src/uart/uart_transmitter.sv