../../src/util/counter.sv