../../src/uart/uart_receiver.sv